module test ();
input a;
endmodule
