module rtl1 ();
endmodule
