module test ();
endmodule
